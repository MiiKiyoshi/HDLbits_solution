//popcount3.v
module top_module( 
    input [2:0] in,
    output [1:0] out );

//0:00, 1:01, 2:10, 3:11
//
//out[0] = 01'2' + 0'12' + 0'1'2 + 012
//       = (01' + 0'1)2' + (0'1' + 01)2  
//
//       = ((0 ^ 1) & ~2) | (~(0 ^ 1) & 2)
//       = 0 ^ 1 ^ 2;
//
//out[1] = 012' + 01'2 + 0'12 + 012
//       = 0(12' + 1'2) + 12
//
//       = 0 & (1 ^ 2) | 1 & 2

assign out[0] = in[0] ^ in[1] ^ in[2];
assign out[1] = in[0] & (in[1] ^ in[2]) | in[1] & in[2];
    
//assign out = in[0] + in[1] + in[2];

endmodule

